�� z     ?��9*@bf@$5�rT�� PCr�\��^v�Zk��^v gATP_1�`���CX�^�i��6� gATP_2�w��%�%_�w�%�%_ aATP_1�x�>A�4!�w�>A�4! aATP_2��S���'������'� bATP_1���w)������w)��� bATP_2��O��y�f�����y�f bATP_3@r�ᰉ�'@sUᰉ�' 2-DPG@o��x���@p�f<t�T 3-DPG@a�a�D@b�a�D PDE